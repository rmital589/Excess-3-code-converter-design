module Inverter(X,XN);

input X;
output XN;

assign XN = ~X;

endmodule
